module ueda

// The start of Ueda.
